module mux32

endmodule