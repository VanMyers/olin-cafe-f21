module bit_counter (in, num)

input wire [7:0] in;
output logic [3:0] num;

logic 